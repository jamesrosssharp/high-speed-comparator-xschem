magic
tech sky130A
magscale 1 2
timestamp 1738141631
<< error_s >>
rect 245 -1527 280 -1493
rect 246 -1546 280 -1527
rect 76 -1905 134 -1899
rect 76 -1939 88 -1905
rect 76 -1945 134 -1939
rect 265 -2041 280 -1546
rect 299 -1580 334 -1546
rect 614 -1580 649 -1546
rect 299 -2041 333 -1580
rect 615 -1599 649 -1580
rect 1001 -1599 1054 -1598
rect 445 -1648 503 -1642
rect 445 -1682 457 -1648
rect 445 -1688 503 -1682
rect 445 -1958 503 -1952
rect 445 -1992 457 -1958
rect 445 -1998 503 -1992
rect 299 -2075 314 -2041
rect 634 -2094 649 -1599
rect 668 -1633 703 -1599
rect 983 -1633 1054 -1599
rect 668 -2094 702 -1633
rect 984 -1634 1054 -1633
rect 1001 -1668 1072 -1634
rect 1352 -1668 1387 -1634
rect 814 -1701 872 -1695
rect 814 -1735 826 -1701
rect 814 -1741 872 -1735
rect 814 -2011 872 -2005
rect 814 -2045 826 -2011
rect 814 -2051 872 -2045
rect 668 -2128 683 -2094
rect 1001 -2147 1071 -1668
rect 1353 -1687 1387 -1668
rect 1183 -1736 1241 -1730
rect 1183 -1770 1195 -1736
rect 1183 -1776 1241 -1770
rect 1183 -2064 1241 -2058
rect 1183 -2098 1195 -2064
rect 1183 -2104 1241 -2098
rect 1001 -2183 1054 -2147
rect 1372 -2200 1387 -1687
rect 1406 -1721 1441 -1687
rect 1721 -1721 1756 -1687
rect 1406 -2200 1440 -1721
rect 1722 -1740 1756 -1721
rect 1552 -1789 1610 -1783
rect 1552 -1823 1564 -1789
rect 1552 -1829 1610 -1823
rect 1552 -2117 1610 -2111
rect 1552 -2151 1564 -2117
rect 1552 -2157 1610 -2151
rect 1406 -2234 1421 -2200
rect 1741 -2253 1756 -1740
rect 1775 -1774 1810 -1740
rect 2090 -1774 2125 -1757
rect 1775 -2253 1809 -1774
rect 2091 -1775 2125 -1774
rect 2091 -1811 2161 -1775
rect 2477 -1811 2530 -1810
rect 1921 -1842 1979 -1836
rect 1921 -1876 1933 -1842
rect 2108 -1845 2179 -1811
rect 2459 -1845 2530 -1811
rect 1921 -1882 1979 -1876
rect 1921 -2170 1979 -2164
rect 1921 -2204 1933 -2170
rect 1921 -2210 1979 -2204
rect 1775 -2287 1790 -2253
rect 2108 -2306 2178 -1845
rect 2460 -1846 2530 -1845
rect 2477 -1880 2548 -1846
rect 2290 -1913 2348 -1907
rect 2290 -1947 2302 -1913
rect 2290 -1953 2348 -1947
rect 2290 -2223 2348 -2217
rect 2290 -2257 2302 -2223
rect 2290 -2263 2348 -2257
rect 2108 -2342 2161 -2306
rect 2477 -2359 2547 -1880
rect 2659 -1948 2717 -1942
rect 2659 -1982 2671 -1948
rect 2659 -1988 2717 -1982
rect 2659 -2276 2717 -2270
rect 2659 -2310 2671 -2276
rect 2659 -2316 2717 -2310
rect 2477 -2395 2530 -2359
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__nfet_01v8_V8CAV6  XM1
timestamp 1738141631
transform 1 0 105 0 1 -1767
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XM2
timestamp 1738141631
transform 1 0 474 0 1 -1820
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XM3
timestamp 1738141631
transform 1 0 843 0 1 -1873
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM4
timestamp 1738141631
transform 1 0 1212 0 1 -1917
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM5
timestamp 1738141631
transform 1 0 1581 0 1 -1970
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM6
timestamp 1738141631
transform 1 0 1950 0 1 -2023
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_V8CAV6  XM7
timestamp 1738141631
transform 1 0 2319 0 1 -2085
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM8
timestamp 1738141631
transform 1 0 2688 0 1 -2129
box -211 -319 211 319
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VLAT_PLUS
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VLAT_MINUS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VOUT
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
