Test bench for high speed comparator

.lib /home/jrsharp/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice sf
.inc /home/jrsharp/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.inc high_speed_comp_top.spice

** Supply voltage
.param VCCGAUSS = agauss(1.8, 0.05, 1)
.param VCC = 'VCCGAUSS'

** Common mode voltage
.param VDLGAUSS = agauss(0.9, 0.33, 1)
.param VDL = VDLGAUSS

** Temperature 
.param TEMPGAUSS = agauss(40, 30, 1)
.option temp = 'TEMPGAUSS'

.param trans_time = agauss(500n, 10n, 1)

.param DELTA = 0.1

E5 TEMPERAT VSS VOL=' temper '

VCLK CLK GND PULSE(0 1.8 0 1NS 1NS 10NS 20NS 0)
VVSS VSS GND 0
VVDD VDD GND 'VCC'

VPLUS INP GND 'VDL'
VMINUS INN GND pwl 0 'VDL-DELTA' 10.5n 'VDL-DELTA' 'trans_time' 'VDL+DELTA' 600n 'VDL+DELTA'

X1 CLK INP INN VDD COMP_OUT VSS high_speed_comp_top 

.control
*  set filetype=ascii 
  setseed  8
  reset
  let run = 1
  save all
  op
  write high_speed_comp_sf.raw
  reset
  set appendwrite
  dowhile run < = 100
    save vdd i(vvdd) temperat clk comp_out inn inp
    *save all
    tran 0.1n 600n uic
    write high_speed_comp_sf.raw
    let run = run + 1
    reset
  end
  quit 0
.endc

