Test bench for ac analysis of RF amp

.lib /home/jrsharp/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ${CORNER}

.inc RF_amp.spice

*.subckt RF_amp VDD VINN VOUT VINP VB VSS
x1 VDD VINN VOUT VINP VB VSS RF_amp  

V1 VDD GND 1.8
VPLUS VINP GND DC 0.9 AC 1
VMINUS VINN GND DC 0.9 AC 0

.param VBGAUSS = unif(0.7, 0.3)
*.param VBGAUSS = 0.85
.param VBIAS = 'VBGAUSS'

V2 VB GND 'VBIAS'
V3 VSS GND 0

.control
  setseed 8
  let run = 1
  op	
  save all
  reset
  set appendwrite
  dowhile run < = 100
    save all
*    save frequency v(vout) v(vb)
    op
    write ${RAW_FILE}
    ac dec 10 1 10G
    write ${RAW_FILE}
    let run = run + 1
    reset
  end
  quit 0

.endc
