magic
tech sky130A
magscale 1 2
timestamp 1738148512
<< error_s >>
rect 1263 -3775 1298 -3741
rect 1264 -3794 1298 -3775
rect 1094 -4153 1152 -4147
rect 1094 -4187 1106 -4153
rect 1094 -4193 1152 -4187
rect 1283 -4289 1298 -3794
rect 1317 -3828 1352 -3794
rect 1632 -3828 1667 -3794
rect 1317 -4289 1351 -3828
rect 1633 -3847 1667 -3828
rect 2019 -3847 2072 -3846
rect 1463 -3896 1521 -3890
rect 1463 -3930 1475 -3896
rect 1463 -3936 1521 -3930
rect 1463 -4206 1521 -4200
rect 1463 -4240 1475 -4206
rect 1463 -4246 1521 -4240
rect 1317 -4323 1332 -4289
rect 1652 -4342 1667 -3847
rect 1686 -3881 1721 -3847
rect 2001 -3881 2072 -3847
rect 1686 -4342 1720 -3881
rect 2002 -3882 2072 -3881
rect 2019 -3916 2090 -3882
rect 2370 -3916 2405 -3882
rect 1832 -3949 1890 -3943
rect 1832 -3983 1844 -3949
rect 1832 -3989 1890 -3983
rect 1832 -4259 1890 -4253
rect 1832 -4293 1844 -4259
rect 1832 -4299 1890 -4293
rect 1686 -4376 1701 -4342
rect 2019 -4395 2089 -3916
rect 2371 -3935 2405 -3916
rect 2201 -3984 2259 -3978
rect 2201 -4018 2213 -3984
rect 2201 -4024 2259 -4018
rect 2201 -4312 2259 -4306
rect 2201 -4346 2213 -4312
rect 2201 -4352 2259 -4346
rect 2019 -4431 2072 -4395
rect 2390 -4448 2405 -3935
rect 2424 -3969 2459 -3935
rect 2739 -3969 2774 -3935
rect 2424 -4448 2458 -3969
rect 2740 -3988 2774 -3969
rect 2570 -4037 2628 -4031
rect 2570 -4071 2582 -4037
rect 2570 -4077 2628 -4071
rect 2570 -4365 2628 -4359
rect 2570 -4399 2582 -4365
rect 2570 -4405 2628 -4399
rect 2424 -4482 2439 -4448
rect 2759 -4501 2774 -3988
rect 2793 -4022 2828 -3988
rect 3108 -4022 3143 -4005
rect 2793 -4501 2827 -4022
rect 3109 -4023 3143 -4022
rect 3109 -4059 3179 -4023
rect 3495 -4059 3548 -4058
rect 2939 -4090 2997 -4084
rect 2939 -4124 2951 -4090
rect 3126 -4093 3197 -4059
rect 3477 -4093 3548 -4059
rect 2939 -4130 2997 -4124
rect 2939 -4418 2997 -4412
rect 2939 -4452 2951 -4418
rect 2939 -4458 2997 -4452
rect 2793 -4535 2808 -4501
rect 3126 -4554 3196 -4093
rect 3478 -4094 3548 -4093
rect 3495 -4128 3566 -4094
rect 3308 -4161 3366 -4155
rect 3308 -4195 3320 -4161
rect 3308 -4201 3366 -4195
rect 3308 -4471 3366 -4465
rect 3308 -4505 3320 -4471
rect 3308 -4511 3366 -4505
rect 3126 -4590 3179 -4554
rect 3495 -4607 3565 -4128
rect 3677 -4196 3735 -4190
rect 3677 -4230 3689 -4196
rect 3677 -4236 3735 -4230
rect 3677 -4524 3735 -4518
rect 3677 -4558 3689 -4524
rect 3677 -4564 3735 -4558
rect 3495 -4643 3548 -4607
rect 3290 -5554 3348 -5548
rect 2870 -5562 2928 -5556
rect 1182 -5576 1240 -5570
rect 1182 -5610 1194 -5576
rect 1604 -5578 1662 -5572
rect 1182 -5616 1240 -5610
rect 1604 -5612 1616 -5578
rect 2870 -5596 2882 -5562
rect 3290 -5588 3302 -5554
rect 3290 -5594 3348 -5588
rect 2870 -5602 2928 -5596
rect 1604 -5618 1662 -5612
rect 2448 -7370 2506 -7364
rect 2026 -7378 2084 -7372
rect 2026 -7412 2038 -7378
rect 2448 -7404 2460 -7370
rect 2448 -7410 2506 -7404
rect 2026 -7418 2084 -7412
rect 3290 -7682 3348 -7676
rect 2870 -7690 2928 -7684
rect 2448 -7698 2506 -7692
rect 1182 -7704 1240 -7698
rect 1182 -7738 1194 -7704
rect 1604 -7706 1662 -7700
rect 2026 -7706 2084 -7700
rect 1182 -7744 1240 -7738
rect 1604 -7740 1616 -7706
rect 2026 -7740 2038 -7706
rect 2448 -7732 2460 -7698
rect 2870 -7724 2882 -7690
rect 3290 -7716 3302 -7682
rect 3290 -7722 3348 -7716
rect 2870 -7730 2928 -7724
rect 2448 -7738 2506 -7732
rect 1604 -7746 1662 -7740
rect 2026 -7746 2084 -7740
rect 2462 -8138 2520 -8132
rect 2030 -8144 2088 -8138
rect 2030 -8178 2042 -8144
rect 2462 -8172 2474 -8138
rect 2462 -8178 2520 -8172
rect 2030 -8184 2088 -8178
rect 2462 -8448 2520 -8442
rect 2030 -8454 2088 -8448
rect 2030 -8488 2042 -8454
rect 2462 -8482 2474 -8448
rect 2462 -8488 2520 -8482
rect 2030 -8494 2088 -8488
<< metal1 >>
rect 1314 -42 1514 158
rect 1748 -24 1948 176
rect 2338 -40 2538 160
rect 4330 26 4530 226
rect 1186 -11452 1386 -11252
rect 1796 -11472 1996 -11272
use strong_arm_latch  x1
timestamp 1738148512
transform 1 0 174 0 1 -6681
box 0 -4381 3356 1265
use post_amplifier  x2
timestamp 1738141631
transform 1 0 1018 0 1 -2248
box -106 -2448 2899 200
use sky130_fd_sc_hd__dfxtp_2  x3 ~/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1738142526
transform 1 0 2704 0 1 -1974
box -38 -48 1602 592
use sky130_fd_sc_hd__clkinv_4  x4 ~/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1728392188
transform 1 0 950 0 1 -1970
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  x5 ~/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1738142205
transform 1 0 1670 0 1 -1970
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  x6 ~/home_mnt/asic/sky130_pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1728392188
transform 1 0 2022 0 1 -1970
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  x7
timestamp 1738142205
transform 1 0 2188 0 1 -1970
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  x8
timestamp 1728392188
transform 1 0 2538 0 1 -1972
box -38 -48 130 592
<< labels >>
flabel metal1 1314 -42 1514 158 0 FreeSans 256 0 0 0 CLK
port 0 nsew
flabel metal1 1748 -24 1948 176 0 FreeSans 256 0 0 0 COMP_OUT
port 4 nsew
flabel metal1 2338 -40 2538 160 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 4330 26 4530 226 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 1186 -11452 1386 -11252 0 FreeSans 256 0 0 0 VINP
port 1 nsew
flabel metal1 1796 -11472 1996 -11272 0 FreeSans 256 0 0 0 VINN
port 2 nsew
<< end >>
