** sch_path: /home/jrsharp/home_mnt/asic/high_speed_comparator/xschem/high_speed_comp_top.sch
.subckt high_speed_comp_top CLK VINP VINN VDD COMP_OUT VSS
*.PININFO VINP:I VINN:I VDD:I VSS:I CLK:I COMP_OUT:O
x1 VDD CLK_PRIME net1 net2 VSS VINP VINN strong_arm_latch
x2 VDD net1 net2 VOUT VSS post_amplifier
x3 CLK VOUT GND GND VDD VDD COMP_OUT sky130_fd_sc_hd__dfxtp_2
x4 CLK GND GND VDD VDD CLK_PRIME sky130_fd_sc_hd__clkinv_4
x5 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
x6 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
x7 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
x8 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
.ends

* expanding   symbol:  strong_arm_latch.sym # of pins=7
** sym_path: /home/jrsharp/home_mnt/asic/high_speed_comparator/xschem/strong_arm_latch.sym
** sch_path: /home/jrsharp/home_mnt/asic/high_speed_comparator/xschem/strong_arm_latch.sch
.subckt strong_arm_latch VDD CLK VOUT_PLUS VOUT_MINUS VSS VINP VINN
*.PININFO VSS:I VDD:I CLK:I VINP:I VINN:I VOUT_MINUS:O VOUT_PLUS:O
XM1 net2 VINP net1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=10 nf=1 m=1
XM2 net3 VINN net1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=10 nf=1 m=1
XM3 net1 CLK VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=10 nf=1 m=1
XM4 VOUT_PLUS VOUT_MINUS net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 VOUT_MINUS VOUT_PLUS net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 VOUT_PLUS VOUT_MINUS VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 VOUT_MINUS VOUT_PLUS VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 VOUT_PLUS CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM9 net2 CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM10 VOUT_MINUS CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
XM11 net3 CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 m=1
.ends


* expanding   symbol:  post_amplifier.sym # of pins=5
** sym_path: /home/jrsharp/home_mnt/asic/high_speed_comparator/xschem/post_amplifier.sym
** sch_path: /home/jrsharp/home_mnt/asic/high_speed_comparator/xschem/post_amplifier.sch
.subckt post_amplifier VDD VLAT_PLUS VLAT_MINUS VOUT VSS
*.PININFO VLAT_PLUS:I VLAT_MINUS:I VDD:I VSS:I VOUT:O
XM1 net1 VLAT_PLUS net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net3 VLAT_MINUS net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net4 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net1 VLAT_PLUS net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net3 VLAT_MINUS net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 VOUT net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 VOUT net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
